package arb_pkg;
    int no_of_trans = 50;
    
    `include "./../env/arb_trans.sv"
    `include "./../env/arb_gen.sv"
    `include "./../env/arb_drv.sv"
    `include "./../env/arb_mon.sv"
    `include "./../env/arb_cov_model.sv"
    `include "./../env/arb_sb.sv"
    `include "./../env/arb_env.sv"
endpackage